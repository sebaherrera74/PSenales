[HEAD]:117
VPP:49639.398438
OFFSET:0.000000
CHANNEL:1
RATEPOS:0.000025
RATENEG:0.000025
MAX:32767.000000
MIN:3147.000000
[DATA]:39
K7[�.!�&�,H28�=�CJI�NET�Y�^Uc�gl�ovs�vQy�{p}�~����}|�y�v)sonj:ez_