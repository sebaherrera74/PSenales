[HEAD]:115
VPP:2.800000
OFFSET:0.000000
CHANNEL:1
RATEPOS:0.000061
RATENEG:0.000061
MAX:32767.000000
MIN:-32767.000000
[DATA]:1000
  X��B|���!�%�)C-�0U4�7�:�=�@lC�EJHgJcL.N�OQ6R,S�StT�T�T�T�TTnS�R�QKP�NHM�K�I�GhE*C�@6>�;�8633G0P-O*I'@$7!22;Ps��Q
�^� ����8���6�������J���s�Q�b�����������]�������� D�f1.]�� "�%{)=-	1�4�8�<Y@1D�G�KeOS�VZ{]�`�c�f�i�l'o�q�s�u�w�y{i|}u~)������~4~>}|�zyZw]uAs�psn�kifc�_�\!Y�URoN�J�FCT?|;�7�3�/0,q(�$!��xQKg
��R 7�G�������^�_������Y�V����x�:�+�K������z�i�|�{	�m="%!(%+$.1 4�6�9S<�>_A�CF)H5JL�MDO�P�Q�R�SCT�T�T�T�TST�S�R�Q�PUO�M�K�I�GGE�B�?=�9�6a3�/=,}(�$� ��Q�y#��t� ����Z�3���7�jպ�)λ�p�L�O����`�#���_�毎�x���ޫk�*��:����Ԭ��Ю���*������+�������*��ǹʛ͋ЅӇ֏٘ܠߤ���}�U����f���I�������=�'Z	`
8�V���>�
��4��� n�����������h���w���5�{ն����:�a�ɺ�;����i�����[�H�F�d���$�ƍ���������E�/�Z���C���3���9���L�Ņ_�:�6�c�A��×Ś؝�`�է[�񮧲^�%�콽���n�D���ԗ�D���g���0�k����a�����G X;�u��	�
�,���e�W�
�	]�� ����M���=��������!�%�!�����	��3�_Ȟ���^�콎�P�D�G�|�ұY�����0���:���[�ͫq�W�]����Ȳ������m��������,ʕ� ��ԓ�v�r�������h����i�]���  �#�'�+G/�236s9�<~?5B�DCG�I�KiMO|P�Q�R�SCT�T�T�T�TST�S�R�Q�P�O�MRL�J�HnF1D�AZ?�<:Q7{4�1�.�+�(�%�"������#x�n�������Q����X�_������Z�U����t�9�0�Y���>�������6�5�	���.��� $$�'�+X/)3�6�:�>vBNFJ�MrQU�X\F_zb�e�h`k n�p�ruw�xlz�{}~�~{����:�~�}�|R{�yxCv6t�q�o�lJjhgfdBa�]�Z5W�S	PRL�H�D�@1=Y9�5�1�-*b&�"$�8�����0�Q"��G���'�������5���j�Q�j��1���������c�������� ��`�	3������ �#�&�)�,�/�2�5g8#;�=I@�BECGPI<KM�N	PQQhRMST�T�T�T�T�TTMShRQQ�OoN�L�J�HNF�C.A^>];48�4s1�-+*[&q"oX/��e	� b����t�7�	��������Zӻ�=��ȬŞ�ȿ�w����$���"����0���:���[�ͫq�F�M����v�1���6�s��\��î�w�R�;�1�0�6�>�G�N�O�G�5�����A���=������ �����	�
�'���i�Z�
�	K�L��o�"����I�a�W�-����
�z���%�dә������?�s����.����}��ԟ�������K�̎��q�u���1�Ƀ������d����d�瀬��������e�Q�m���*���{�m�o����L���W�����k�B��