[HEAD]:115
VPP:2.800000
OFFSET:0.000000
CHANNEL:1
RATEPOS:0.000059
RATENEG:0.000059
MAX:18863.000000
MIN:-32768.000000
[DATA]:1000
�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A            �A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$���I� � �I�����$�A�I�>I(����I(�>�I�A�$