[HEAD]:115
VPP:2.800000
OFFSET:0.000000
CHANNEL:1
RATEPOS:0.000061
RATENEG:0.000061
MAX:32767.000000
MIN:-32767.000000
[DATA]:500
�%�����D�m���G��)3=OP�aKp�z���zKp�aOP3=�)�G��m�D�������%�4iB�L�SDU�QI�; *�  3���e��6���y�	����-�e�H�|�	��
m��B�*��±�0���i���i���0�����*�B��m�
��	|H�e�-�˗�	�y���6��e���3�              �%�����D�m���G��)3=OP�aKp�z���zKp�aOP3=�)�G��m�D�������%�4iB�L�SDU�QI�; *�  3���e��6���y�	����-�e�H�|�	��
m��B�*��±�0���i���i���0�����*�B��m�
��	|H�e�-�˗�	�y���6��e���3�              �%�����D�m���G��)3=OP�aKp�z���zKp�aOP3=�)�G��m�D�������%�4iB�L�SDU�QI�; *�  3���e��6���y�	����-�e�H�|�	��
m��B�*��±�0���i���i���0�����*�B��m�
��	|H�e�-�˗�	�y���6��e���3�              �%�����D�m���G��)3=OP�aKp�z���zKp�aOP3=�)�G��m�D�������%�4iB�L�SDU�QI�; *�  3���e��6���y�	����-�e�H�|�	��
m��B�*��±�0���i���i���0�����*�B��m�
��	|H�e�-�˗�	�y���6��e���3�              �%�����D�m���G��)3=OP�aKp�z���zKp�aOP3=�)�G��m�D�������%�4iB�L�SDU�QI�; *�  3���e��6���y�	����-�e�H�|�	��
m��B�*��±�0���i���i���0�